// *****************************************************
// AVR address constants (localparams)
//  for registers used by Xcelerator Blocks (XBs) 
// *****************************************************

localparam SVCR_ADDR  = 8'hFA;
localparam SVPWL_ADDR = 8'hFC;
localparam SVPWH_ADDR = 8'hFD;

